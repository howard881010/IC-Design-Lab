module Alpha_table(
input clk,
input srstn,
input [7:0] alpha_a,
input [7:0] alpha_b,
input [7:0] alpha_c,
input [7:0] alpha_d,
input [7:0] value_e,
input [7:0] value_f,
input [7:0] value_g,
input [7:0] value_h,
input [7:0] alpha_i,
//input err_correct_en,

output reg [7:0] value_a,
output reg [7:0] value_b,
output reg [7:0] value_c,
output reg [7:0] value_d,
output reg [7:0] alpha_e,
output reg [7:0] alpha_f,
output reg [7:0] alpha_g,
output reg [7:0] alpha_h,
output reg [7:0] value_i
///output reg find_done
);

reg [7:0] new_value_a, new_value_b, new_value_c, new_value_d, new_alpha_e, new_alpha_f, new_alpha_g, new_alpha_h, new_value_i;

always @(posedge clk) begin
	if(~srstn) begin
        value_a <= 0;
        value_b <= 0;
        value_c <= 0;
        value_d <= 0;
        alpha_e <= 0;
        alpha_f <= 0;
        alpha_g <= 0;
        alpha_h <= 0;
        value_i <= 0;

    end
    else begin 
        
        value_a <= new_value_a;
        value_b <= new_value_b;
        value_c <= new_value_c;
        value_d <= new_value_d;
        //if (new_alpha_e != 0)
            alpha_e <= new_alpha_e;
        //else 
           // alpha_e <= alpha_e;
        //if (new_alpha_f != 0)
            alpha_f <= new_alpha_f;
        //else 
            //alpha_f <= alpha_f;
       // if(new_alpha_g != 0)
            alpha_g <= new_alpha_g;
        //else 
           // alpha_g <= alpha_g;
       // if (new_alpha_h != 0)
            alpha_h <= new_alpha_h;
        //else    
           // alpha_h <= alpha_h;
           value_i <= new_value_i;
    end
end

always @* begin
    case(alpha_a) //synopsys parallel_case
        0: new_value_a =  1;
        1: new_value_a =  2;
        2: new_value_a =  4;
        3: new_value_a =  8;
        4: new_value_a =  16;
        5: new_value_a =  32;
        6: new_value_a =  64;
        7: new_value_a =  128;
        8: new_value_a =  29;
        9: new_value_a =  58;
        10: new_value_a =  116;
        11: new_value_a =  232;
        12: new_value_a =  205;
        13: new_value_a =  135;
        14: new_value_a =  19;
        15: new_value_a =  38;
        16: new_value_a =  76;
        17: new_value_a =  152;
        18: new_value_a =  45;
        19: new_value_a =  90;
        20: new_value_a =  180;
        21: new_value_a =  117;
        22: new_value_a = 	234;
        23: new_value_a = 	201;
        24: new_value_a = 	143;
        25: new_value_a = 	3;
        26: new_value_a = 	6;
        27: new_value_a = 	12;
        28: new_value_a = 	24;
        29: new_value_a = 	48;
        30: new_value_a = 	96;
        31: new_value_a = 	192;
        32: new_value_a = 	157;
        33: new_value_a = 	39;
        34: new_value_a = 	78;
        35: new_value_a = 	156;
        36: new_value_a = 	37;
        37: new_value_a = 	74;
        38: new_value_a = 	148;
        39: new_value_a = 	53;
        40: new_value_a = 	106;
        41: new_value_a = 	212;
        42: new_value_a = 	181;
        43: new_value_a = 	119;
        44: new_value_a = 	238;
        45: new_value_a = 	193;
        46: new_value_a = 	159;
        47: new_value_a = 	35;
        48: new_value_a = 	70;
        49: new_value_a = 	140;
        50: new_value_a = 	5;
        51: new_value_a = 	10;
        52: new_value_a = 	20;
        53: new_value_a = 	40;
        54: new_value_a = 	80;
        55: new_value_a = 	160;
        56: new_value_a = 	93;
        57: new_value_a = 	186;
        58: new_value_a = 	105;
        59: new_value_a = 	210;
        60: new_value_a = 	185;
        61: new_value_a = 	111;
        62: new_value_a = 	222;
        63: new_value_a = 	161;
        64: new_value_a = 	95;
        65: new_value_a = 	190;
        66: new_value_a = 	97;
        67: new_value_a = 	194;
        68: new_value_a = 	153;
        69: new_value_a = 	47;
        70: new_value_a = 	94;
        71: new_value_a = 	188;
        72: new_value_a = 	101;
        73: new_value_a = 	202;
        74: new_value_a = 	137;
        75: new_value_a = 	15;
        76: new_value_a = 	30;
        77: new_value_a = 	60;
        78: new_value_a = 	120;
        79: new_value_a = 	240;
        80: new_value_a = 	253;
        81: new_value_a = 	231;
        82: new_value_a = 	211;
        83: new_value_a = 	187;
        84: new_value_a = 	107;
        85: new_value_a = 	214;
        86: new_value_a = 	177;
        87: new_value_a = 	127;
        88: new_value_a = 	254;
        89: new_value_a = 	225;
        90: new_value_a = 	223;
        91: new_value_a = 	163;
        92: new_value_a = 	91;
        93: new_value_a = 	182;
        94: new_value_a = 	113;
        95: new_value_a = 	226;
        96: new_value_a = 	217;
        97: new_value_a = 	175;
        98: new_value_a = 	67;
        99: new_value_a = 	134;
        100: new_value_a = 	17;
        101: new_value_a = 	34;
        102: new_value_a = 	68;
        103: new_value_a = 	136;
        104: new_value_a = 	13;
        105: new_value_a = 	26;
        106: new_value_a = 	52;
        107: new_value_a = 	104;
        108: new_value_a = 	208;
        109: new_value_a = 	189;
        110: new_value_a = 	103;
        111: new_value_a = 	206;
        112: new_value_a = 	129;
        113: new_value_a = 	31;
        114: new_value_a = 	62;
        115: new_value_a = 	124;
        116: new_value_a = 	248;
        117: new_value_a = 	237;
        118: new_value_a = 	199;
        119: new_value_a = 	147;
        120: new_value_a = 	59;
        121: new_value_a = 	118;
        122: new_value_a = 	236;
        123: new_value_a = 	197;
        124: new_value_a = 	151;
        125: new_value_a = 	51;
        126: new_value_a = 	102;
        127: new_value_a = 	204;
        128: new_value_a = 	133;
        129: new_value_a = 	23;
        130: new_value_a = 	46;
        131: new_value_a = 	92;
        132: new_value_a = 	184;
        133: new_value_a = 	109;
        134: new_value_a = 	218;
        135: new_value_a = 	169;
        136: new_value_a = 	79;
        137: new_value_a = 	158;
        138: new_value_a = 	33;
        139: new_value_a = 	66;
        140: new_value_a = 	132;
        141: new_value_a = 	21;
        142: new_value_a = 	42;
        143: new_value_a = 	84;
        144: new_value_a = 	168;
        145: new_value_a = 	77;
        146: new_value_a = 	154;
        147: new_value_a = 	41;
        148: new_value_a = 	82;
        149: new_value_a = 	164;
        150: new_value_a = 	85;
        151: new_value_a = 	170;
        152: new_value_a = 	73;
        153: new_value_a = 	146;
        154: new_value_a = 	57;
        155: new_value_a = 	114;
        156: new_value_a = 	228;
        157: new_value_a = 	213;
        158: new_value_a = 	183;
        159: new_value_a = 	115;
        160: new_value_a = 	230;
        161: new_value_a = 	209;
        162: new_value_a = 	191;
        163: new_value_a = 	99;
        164: new_value_a = 	198;
        165: new_value_a = 	145;
        166: new_value_a = 	63;
        167: new_value_a = 	126;
        168: new_value_a = 	252;
        169: new_value_a = 	229;
        170: new_value_a = 	215;
        171: new_value_a = 	179;
        172: new_value_a = 	123;
        173: new_value_a = 	246;
        174: new_value_a = 	241;
        175: new_value_a = 	255;
        176: new_value_a = 	227;
        177: new_value_a = 	219;
        178: new_value_a = 	171;
        179: new_value_a = 	75;
        180: new_value_a = 	150;
        181: new_value_a = 	49;
        182: new_value_a = 	98;
        183: new_value_a = 	196;
        184: new_value_a = 	149;
        185: new_value_a = 	55;
        186: new_value_a = 	110;
        187: new_value_a = 	220;
        188: new_value_a = 	165;
        189: new_value_a = 	87;
        190: new_value_a = 	174;
        191: new_value_a = 	65;
        192: new_value_a = 	130;
        193: new_value_a = 	25;
        194: new_value_a = 	50;
        195: new_value_a = 	100;
        196: new_value_a = 	200;
        197: new_value_a = 	141;
        198: new_value_a = 	7;
        199: new_value_a = 	14;
        200: new_value_a = 	28;
        201: new_value_a = 	56;
        202: new_value_a = 	112;
        203: new_value_a = 	224;
        204: new_value_a = 	221;
        205: new_value_a = 	167;
        206: new_value_a = 	83;
        207: new_value_a = 	166;
        208: new_value_a = 	81;
        209: new_value_a = 	162;
        210: new_value_a = 	89;
        211: new_value_a = 	178;
        212: new_value_a = 	121;
        213: new_value_a = 	242;
        214: new_value_a = 	249;
        215: new_value_a = 	239;
        216: new_value_a = 	195;
        217: new_value_a = 	155;
        218: new_value_a = 	43;
        219: new_value_a = 	86;
        220: new_value_a = 	172;
        221: new_value_a = 	69;
        222: new_value_a = 	138;
        223: new_value_a = 	9;
        224: new_value_a = 	18;
        225: new_value_a = 	36;
        226: new_value_a = 	72;
        227: new_value_a = 	144;
        228: new_value_a = 	61;
        229: new_value_a = 	122;
        230: new_value_a = 	244;
        231: new_value_a = 	245;
        232: new_value_a = 	247;
        233: new_value_a = 	243;
        234: new_value_a = 	251;
        235: new_value_a = 	235;
        236: new_value_a = 	203;
        237: new_value_a = 	139;
        238: new_value_a = 	11;
        239: new_value_a = 	22;
        240: new_value_a = 	44;
        241: new_value_a = 	88;
        242: new_value_a = 	176;
        243: new_value_a = 	125;
        244: new_value_a = 	250;
        245: new_value_a = 	233;
        246: new_value_a = 	207;
        247: new_value_a = 	131;
        248: new_value_a = 	27;
        249: new_value_a = 	54;
        250: new_value_a = 	108;
        251: new_value_a = 	216;
        252: new_value_a = 	173;
        253: new_value_a = 	71;
        254: new_value_a = 	142;
        default: new_value_a = 0;
    endcase
end

always @* begin
    case(alpha_i) //synopsys parallel_case
        0: new_value_i =  1;
        1: new_value_i =  2;
        2: new_value_i =  4;
        3: new_value_i =  8;
        4: new_value_i =  16;
        5: new_value_i =  32;
        6: new_value_i =  64;
        7: new_value_i =  128;
        8: new_value_i =  29;
        9: new_value_i =  58;
        10: new_value_i =  116;
        11: new_value_i =  232;
        12: new_value_i =  205;
        13: new_value_i =  135;
        14: new_value_i =  19;
        15: new_value_i =  38;
        16: new_value_i =  76;
        17: new_value_i =  152;
        18: new_value_i =  45;
        19: new_value_i =  90;
        20: new_value_i =  180;
        21: new_value_i =  117;
        22: new_value_i = 	234;
        23: new_value_i = 	201;
        24: new_value_i = 	143;
        25: new_value_i = 	3;
        26: new_value_i = 	6;
        27: new_value_i = 	12;
        28: new_value_i = 	24;
        29: new_value_i = 	48;
        30: new_value_i = 	96;
        31: new_value_i = 	192;
        32: new_value_i = 	157;
        33: new_value_i = 	39;
        34: new_value_i = 	78;
        35: new_value_i = 	156;
        36: new_value_i = 	37;
        37: new_value_i = 	74;
        38: new_value_i = 	148;
        39: new_value_i = 	53;
        40: new_value_i = 	106;
        41: new_value_i = 	212;
        42: new_value_i = 	181;
        43: new_value_i = 	119;
        44: new_value_i = 	238;
        45: new_value_i = 	193;
        46: new_value_i = 	159;
        47: new_value_i = 	35;
        48: new_value_i = 	70;
        49: new_value_i = 	140;
        50: new_value_i = 	5;
        51: new_value_i = 	10;
        52: new_value_i = 	20;
        53: new_value_i = 	40;
        54: new_value_i = 	80;
        55: new_value_i = 	160;
        56: new_value_i = 	93;
        57: new_value_i = 	186;
        58: new_value_i = 	105;
        59: new_value_i = 	210;
        60: new_value_i = 	185;
        61: new_value_i = 	111;
        62: new_value_i = 	222;
        63: new_value_i = 	161;
        64: new_value_i = 	95;
        65: new_value_i = 	190;
        66: new_value_i = 	97;
        67: new_value_i = 	194;
        68: new_value_i = 	153;
        69: new_value_i = 	47;
        70: new_value_i = 	94;
        71: new_value_i = 	188;
        72: new_value_i = 	101;
        73: new_value_i = 	202;
        74: new_value_i = 	137;
        75: new_value_i = 	15;
        76: new_value_i = 	30;
        77: new_value_i = 	60;
        78: new_value_i = 	120;
        79: new_value_i = 	240;
        80: new_value_i = 	253;
        81: new_value_i = 	231;
        82: new_value_i = 	211;
        83: new_value_i = 	187;
        84: new_value_i = 	107;
        85: new_value_i = 	214;
        86: new_value_i = 	177;
        87: new_value_i = 	127;
        88: new_value_i = 	254;
        89: new_value_i = 	225;
        90: new_value_i = 	223;
        91: new_value_i = 	163;
        92: new_value_i = 	91;
        93: new_value_i = 	182;
        94: new_value_i = 	113;
        95: new_value_i = 	226;
        96: new_value_i = 	217;
        97: new_value_i = 	175;
        98: new_value_i = 	67;
        99: new_value_i = 	134;
        100: new_value_i = 	17;
        101: new_value_i = 	34;
        102: new_value_i = 	68;
        103: new_value_i = 	136;
        104: new_value_i = 	13;
        105: new_value_i = 	26;
        106: new_value_i = 	52;
        107: new_value_i = 	104;
        108: new_value_i = 	208;
        109: new_value_i = 	189;
        110: new_value_i = 	103;
        111: new_value_i = 	206;
        112: new_value_i = 	129;
        113: new_value_i = 	31;
        114: new_value_i = 	62;
        115: new_value_i = 	124;
        116: new_value_i = 	248;
        117: new_value_i = 	237;
        118: new_value_i = 	199;
        119: new_value_i = 	147;
        120: new_value_i = 	59;
        121: new_value_i = 	118;
        122: new_value_i = 	236;
        123: new_value_i = 	197;
        124: new_value_i = 	151;
        125: new_value_i = 	51;
        126: new_value_i = 	102;
        127: new_value_i = 	204;
        128: new_value_i = 	133;
        129: new_value_i = 	23;
        130: new_value_i = 	46;
        131: new_value_i = 	92;
        132: new_value_i = 	184;
        133: new_value_i = 	109;
        134: new_value_i = 	218;
        135: new_value_i = 	169;
        136: new_value_i = 	79;
        137: new_value_i = 	158;
        138: new_value_i = 	33;
        139: new_value_i = 	66;
        140: new_value_i = 	132;
        141: new_value_i = 	21;
        142: new_value_i = 	42;
        143: new_value_i = 	84;
        144: new_value_i = 	168;
        145: new_value_i = 	77;
        146: new_value_i = 	154;
        147: new_value_i = 	41;
        148: new_value_i = 	82;
        149: new_value_i = 	164;
        150: new_value_i = 	85;
        151: new_value_i = 	170;
        152: new_value_i = 	73;
        153: new_value_i = 	146;
        154: new_value_i = 	57;
        155: new_value_i = 	114;
        156: new_value_i = 	228;
        157: new_value_i = 	213;
        158: new_value_i = 	183;
        159: new_value_i = 	115;
        160: new_value_i = 	230;
        161: new_value_i = 	209;
        162: new_value_i = 	191;
        163: new_value_i = 	99;
        164: new_value_i = 	198;
        165: new_value_i = 	145;
        166: new_value_i = 	63;
        167: new_value_i = 	126;
        168: new_value_i = 	252;
        169: new_value_i = 	229;
        170: new_value_i = 	215;
        171: new_value_i = 	179;
        172: new_value_i = 	123;
        173: new_value_i = 	246;
        174: new_value_i = 	241;
        175: new_value_i = 	255;
        176: new_value_i = 	227;
        177: new_value_i = 	219;
        178: new_value_i = 	171;
        179: new_value_i = 	75;
        180: new_value_i = 	150;
        181: new_value_i = 	49;
        182: new_value_i = 	98;
        183: new_value_i = 	196;
        184: new_value_i = 	149;
        185: new_value_i = 	55;
        186: new_value_i = 	110;
        187: new_value_i = 	220;
        188: new_value_i = 	165;
        189: new_value_i = 	87;
        190: new_value_i = 	174;
        191: new_value_i = 	65;
        192: new_value_i = 	130;
        193: new_value_i = 	25;
        194: new_value_i = 	50;
        195: new_value_i = 	100;
        196: new_value_i = 	200;
        197: new_value_i = 	141;
        198: new_value_i = 	7;
        199: new_value_i = 	14;
        200: new_value_i = 	28;
        201: new_value_i = 	56;
        202: new_value_i = 	112;
        203: new_value_i = 	224;
        204: new_value_i = 	221;
        205: new_value_i = 	167;
        206: new_value_i = 	83;
        207: new_value_i = 	166;
        208: new_value_i = 	81;
        209: new_value_i = 	162;
        210: new_value_i = 	89;
        211: new_value_i = 	178;
        212: new_value_i = 	121;
        213: new_value_i = 	242;
        214: new_value_i = 	249;
        215: new_value_i = 	239;
        216: new_value_i = 	195;
        217: new_value_i = 	155;
        218: new_value_i = 	43;
        219: new_value_i = 	86;
        220: new_value_i = 	172;
        221: new_value_i = 	69;
        222: new_value_i = 	138;
        223: new_value_i = 	9;
        224: new_value_i = 	18;
        225: new_value_i = 	36;
        226: new_value_i = 	72;
        227: new_value_i = 	144;
        228: new_value_i = 	61;
        229: new_value_i = 	122;
        230: new_value_i = 	244;
        231: new_value_i = 	245;
        232: new_value_i = 	247;
        233: new_value_i = 	243;
        234: new_value_i = 	251;
        235: new_value_i = 	235;
        236: new_value_i = 	203;
        237: new_value_i = 	139;
        238: new_value_i = 	11;
        239: new_value_i = 	22;
        240: new_value_i = 	44;
        241: new_value_i = 	88;
        242: new_value_i = 	176;
        243: new_value_i = 	125;
        244: new_value_i = 	250;
        245: new_value_i = 	233;
        246: new_value_i = 	207;
        247: new_value_i = 	131;
        248: new_value_i = 	27;
        249: new_value_i = 	54;
        250: new_value_i = 	108;
        251: new_value_i = 	216;
        252: new_value_i = 	173;
        253: new_value_i = 	71;
        254: new_value_i = 	142;
        default: new_value_i = 0;
    endcase
end

always @* begin
    case(alpha_b) //synopsys parallel_case
        0: new_value_b =  1;
        1: new_value_b =  2;
        2: new_value_b =  4;
        3: new_value_b =  8;
        4: new_value_b =  16;
        5: new_value_b =  32;
        6: new_value_b =  64;
        7: new_value_b =  128;
        8: new_value_b =  29;
        9: new_value_b =  58;
        10: new_value_b =  116;
        11: new_value_b =  232;
        12: new_value_b =  205;
        13: new_value_b =  135;
        14: new_value_b =  19;
        15: new_value_b =  38;
        16: new_value_b =  76;
        17: new_value_b =  152;
        18: new_value_b =  45;
        19: new_value_b =  90;
        20: new_value_b =  180;
        21: new_value_b =  117;
        22: new_value_b = 	234;
        23: new_value_b = 	201;
        24: new_value_b = 	143;
        25: new_value_b = 	3;
        26: new_value_b = 	6;
        27: new_value_b = 	12;
        28: new_value_b = 	24;
        29: new_value_b = 	48;
        30: new_value_b = 	96;
        31: new_value_b = 	192;
        32: new_value_b = 	157;
        33: new_value_b = 	39;
        34: new_value_b = 	78;
        35: new_value_b = 	156;
        36: new_value_b = 	37;
        37: new_value_b = 	74;
        38: new_value_b = 	148;
        39: new_value_b = 	53;
        40: new_value_b = 	106;
        41: new_value_b = 	212;
        42: new_value_b = 	181;
        43: new_value_b = 	119;
        44: new_value_b = 	238;
        45: new_value_b = 	193;
        46: new_value_b = 	159;
        47: new_value_b = 	35;
        48: new_value_b = 	70;
        49: new_value_b = 	140;
        50: new_value_b = 	5;
        51: new_value_b = 	10;
        52: new_value_b = 	20;
        53: new_value_b = 	40;
        54: new_value_b = 	80;
        55: new_value_b = 	160;
        56: new_value_b = 	93;
        57: new_value_b = 	186;
        58: new_value_b = 	105;
        59: new_value_b = 	210;
        60: new_value_b = 	185;
        61: new_value_b = 	111;
        62: new_value_b = 	222;
        63: new_value_b = 	161;
        64: new_value_b = 	95;
        65: new_value_b = 	190;
        66: new_value_b = 	97;
        67: new_value_b = 	194;
        68: new_value_b = 	153;
        69: new_value_b = 	47;
        70: new_value_b = 	94;
        71: new_value_b = 	188;
        72: new_value_b = 	101;
        73: new_value_b = 	202;
        74: new_value_b = 	137;
        75: new_value_b = 	15;
        76: new_value_b = 	30;
        77: new_value_b = 	60;
        78: new_value_b = 	120;
        79: new_value_b = 	240;
        80: new_value_b = 	253;
        81: new_value_b = 	231;
        82: new_value_b = 	211;
        83: new_value_b = 	187;
        84: new_value_b = 	107;
        85: new_value_b = 	214;
        86: new_value_b = 	177;
        87: new_value_b = 	127;
        88: new_value_b = 	254;
        89: new_value_b = 	225;
        90: new_value_b = 	223;
        91: new_value_b = 	163;
        92: new_value_b = 	91;
        93: new_value_b = 	182;
        94: new_value_b = 	113;
        95: new_value_b = 	226;
        96: new_value_b = 	217;
        97: new_value_b = 	175;
        98: new_value_b = 	67;
        99: new_value_b = 	134;
        100: new_value_b = 	17;
        101: new_value_b = 	34;
        102: new_value_b = 	68;
        103: new_value_b = 	136;
        104: new_value_b = 	13;
        105: new_value_b = 	26;
        106: new_value_b = 	52;
        107: new_value_b = 	104;
        108: new_value_b = 	208;
        109: new_value_b = 	189;
        110: new_value_b = 	103;
        111: new_value_b = 	206;
        112: new_value_b = 	129;
        113: new_value_b = 	31;
        114: new_value_b = 	62;
        115: new_value_b = 	124;
        116: new_value_b = 	248;
        117: new_value_b = 	237;
        118: new_value_b = 	199;
        119: new_value_b = 	147;
        120: new_value_b = 	59;
        121: new_value_b = 	118;
        122: new_value_b = 	236;
        123: new_value_b = 	197;
        124: new_value_b = 	151;
        125: new_value_b = 	51;
        126: new_value_b = 	102;
        127: new_value_b = 	204;
        128: new_value_b = 	133;
        129: new_value_b = 	23;
        130: new_value_b = 	46;
        131: new_value_b = 	92;
        132: new_value_b = 	184;
        133: new_value_b = 	109;
        134: new_value_b = 	218;
        135: new_value_b = 	169;
        136: new_value_b = 	79;
        137: new_value_b = 	158;
        138: new_value_b = 	33;
        139: new_value_b = 	66;
        140: new_value_b = 	132;
        141: new_value_b = 	21;
        142: new_value_b = 	42;
        143: new_value_b = 	84;
        144: new_value_b = 	168;
        145: new_value_b = 	77;
        146: new_value_b = 	154;
        147: new_value_b = 	41;
        148: new_value_b = 	82;
        149: new_value_b = 	164;
        150: new_value_b = 	85;
        151: new_value_b = 	170;
        152: new_value_b = 	73;
        153: new_value_b = 	146;
        154: new_value_b = 	57;
        155: new_value_b = 	114;
        156: new_value_b = 	228;
        157: new_value_b = 	213;
        158: new_value_b = 	183;
        159: new_value_b = 	115;
        160: new_value_b = 	230;
        161: new_value_b = 	209;
        162: new_value_b = 	191;
        163: new_value_b = 	99;
        164: new_value_b = 	198;
        165: new_value_b = 	145;
        166: new_value_b = 	63;
        167: new_value_b = 	126;
        168: new_value_b = 	252;
        169: new_value_b = 	229;
        170: new_value_b = 	215;
        171: new_value_b = 	179;
        172: new_value_b = 	123;
        173: new_value_b = 	246;
        174: new_value_b = 	241;
        175: new_value_b = 	255;
        176: new_value_b = 	227;
        177: new_value_b = 	219;
        178: new_value_b = 	171;
        179: new_value_b = 	75;
        180: new_value_b = 	150;
        181: new_value_b = 	49;
        182: new_value_b = 	98;
        183: new_value_b = 	196;
        184: new_value_b = 	149;
        185: new_value_b = 	55;
        186: new_value_b = 	110;
        187: new_value_b = 	220;
        188: new_value_b = 	165;
        189: new_value_b = 	87;
        190: new_value_b = 	174;
        191: new_value_b = 	65;
        192: new_value_b = 	130;
        193: new_value_b = 	25;
        194: new_value_b = 	50;
        195: new_value_b = 	100;
        196: new_value_b = 	200;
        197: new_value_b = 	141;
        198: new_value_b = 	7;
        199: new_value_b = 	14;
        200: new_value_b = 	28;
        201: new_value_b = 	56;
        202: new_value_b = 	112;
        203: new_value_b = 	224;
        204: new_value_b = 	221;
        205: new_value_b = 	167;
        206: new_value_b = 	83;
        207: new_value_b = 	166;
        208: new_value_b = 	81;
        209: new_value_b = 	162;
        210: new_value_b = 	89;
        211: new_value_b = 	178;
        212: new_value_b = 	121;
        213: new_value_b = 	242;
        214: new_value_b = 	249;
        215: new_value_b = 	239;
        216: new_value_b = 	195;
        217: new_value_b = 	155;
        218: new_value_b = 	43;
        219: new_value_b = 	86;
        220: new_value_b = 	172;
        221: new_value_b = 	69;
        222: new_value_b = 	138;
        223: new_value_b = 	9;
        224: new_value_b = 	18;
        225: new_value_b = 	36;
        226: new_value_b = 	72;
        227: new_value_b = 	144;
        228: new_value_b = 	61;
        229: new_value_b = 	122;
        230: new_value_b = 	244;
        231: new_value_b = 	245;
        232: new_value_b = 	247;
        233: new_value_b = 	243;
        234: new_value_b = 	251;
        235: new_value_b = 	235;
        236: new_value_b = 	203;
        237: new_value_b = 	139;
        238: new_value_b = 	11;
        239: new_value_b = 	22;
        240: new_value_b = 	44;
        241: new_value_b = 	88;
        242: new_value_b = 	176;
        243: new_value_b = 	125;
        244: new_value_b = 	250;
        245: new_value_b = 	233;
        246: new_value_b = 	207;
        247: new_value_b = 	131;
        248: new_value_b = 	27;
        249: new_value_b = 	54;
        250: new_value_b = 	108;
        251: new_value_b = 	216;
        252: new_value_b = 	173;
        253: new_value_b = 	71;
        254: new_value_b = 	142;
        default: new_value_b = 0;
    endcase
end

always @* begin
    case(alpha_c) //synopsys parallel_case
        0: new_value_c =  1;
        1: new_value_c =  2;
        2: new_value_c =  4;
        3: new_value_c =  8;
        4: new_value_c =  16;
        5: new_value_c =  32;
        6: new_value_c =  64;
        7: new_value_c =  128;
        8: new_value_c =  29;
        9: new_value_c =  58;
        10: new_value_c =  116;
        11: new_value_c =  232;
        12: new_value_c =  205;
        13: new_value_c =  135;
        14: new_value_c =  19;
        15: new_value_c =  38;
        16: new_value_c =  76;
        17: new_value_c =  152;
        18: new_value_c =  45;
        19: new_value_c =  90;
        20: new_value_c =  180;
        21: new_value_c =  117;
        22: new_value_c = 	234;
        23: new_value_c = 	201;
        24: new_value_c = 	143;
        25: new_value_c = 	3;
        26: new_value_c = 	6;
        27: new_value_c = 	12;
        28: new_value_c = 	24;
        29: new_value_c = 	48;
        30: new_value_c = 	96;
        31: new_value_c = 	192;
        32: new_value_c = 	157;
        33: new_value_c = 	39;
        34: new_value_c = 	78;
        35: new_value_c = 	156;
        36: new_value_c = 	37;
        37: new_value_c = 	74;
        38: new_value_c = 	148;
        39: new_value_c = 	53;
        40: new_value_c = 	106;
        41: new_value_c = 	212;
        42: new_value_c = 	181;
        43: new_value_c = 	119;
        44: new_value_c = 	238;
        45: new_value_c = 	193;
        46: new_value_c = 	159;
        47: new_value_c = 	35;
        48: new_value_c = 	70;
        49: new_value_c = 	140;
        50: new_value_c = 	5;
        51: new_value_c = 	10;
        52: new_value_c = 	20;
        53: new_value_c = 	40;
        54: new_value_c = 	80;
        55: new_value_c = 	160;
        56: new_value_c = 	93;
        57: new_value_c = 	186;
        58: new_value_c = 	105;
        59: new_value_c = 	210;
        60: new_value_c = 	185;
        61: new_value_c = 	111;
        62: new_value_c = 	222;
        63: new_value_c = 	161;
        64: new_value_c = 	95;
        65: new_value_c = 	190;
        66: new_value_c = 	97;
        67: new_value_c = 	194;
        68: new_value_c = 	153;
        69: new_value_c = 	47;
        70: new_value_c = 	94;
        71: new_value_c = 	188;
        72: new_value_c = 	101;
        73: new_value_c = 	202;
        74: new_value_c = 	137;
        75: new_value_c = 	15;
        76: new_value_c = 	30;
        77: new_value_c = 	60;
        78: new_value_c = 	120;
        79: new_value_c = 	240;
        80: new_value_c = 	253;
        81: new_value_c = 	231;
        82: new_value_c = 	211;
        83: new_value_c = 	187;
        84: new_value_c = 	107;
        85: new_value_c = 	214;
        86: new_value_c = 	177;
        87: new_value_c = 	127;
        88: new_value_c = 	254;
        89: new_value_c = 	225;
        90: new_value_c = 	223;
        91: new_value_c = 	163;
        92: new_value_c = 	91;
        93: new_value_c = 	182;
        94: new_value_c = 	113;
        95: new_value_c = 	226;
        96: new_value_c = 	217;
        97: new_value_c = 	175;
        98: new_value_c = 	67;
        99: new_value_c = 	134;
        100: new_value_c = 	17;
        101: new_value_c = 	34;
        102: new_value_c = 	68;
        103: new_value_c = 	136;
        104: new_value_c = 	13;
        105: new_value_c = 	26;
        106: new_value_c = 	52;
        107: new_value_c = 	104;
        108: new_value_c = 	208;
        109: new_value_c = 	189;
        110: new_value_c = 	103;
        111: new_value_c = 	206;
        112: new_value_c = 	129;
        113: new_value_c = 	31;
        114: new_value_c = 	62;
        115: new_value_c = 	124;
        116: new_value_c = 	248;
        117: new_value_c = 	237;
        118: new_value_c = 	199;
        119: new_value_c = 	147;
        120: new_value_c = 	59;
        121: new_value_c = 	118;
        122: new_value_c = 	236;
        123: new_value_c = 	197;
        124: new_value_c = 	151;
        125: new_value_c = 	51;
        126: new_value_c = 	102;
        127: new_value_c = 	204;
        128: new_value_c = 	133;
        129: new_value_c = 	23;
        130: new_value_c = 	46;
        131: new_value_c = 	92;
        132: new_value_c = 	184;
        133: new_value_c = 	109;
        134: new_value_c = 	218;
        135: new_value_c = 	169;
        136: new_value_c = 	79;
        137: new_value_c = 	158;
        138: new_value_c = 	33;
        139: new_value_c = 	66;
        140: new_value_c = 	132;
        141: new_value_c = 	21;
        142: new_value_c = 	42;
        143: new_value_c = 	84;
        144: new_value_c = 	168;
        145: new_value_c = 	77;
        146: new_value_c = 	154;
        147: new_value_c = 	41;
        148: new_value_c = 	82;
        149: new_value_c = 	164;
        150: new_value_c = 	85;
        151: new_value_c = 	170;
        152: new_value_c = 	73;
        153: new_value_c = 	146;
        154: new_value_c = 	57;
        155: new_value_c = 	114;
        156: new_value_c = 	228;
        157: new_value_c = 	213;
        158: new_value_c = 	183;
        159: new_value_c = 	115;
        160: new_value_c = 	230;
        161: new_value_c = 	209;
        162: new_value_c = 	191;
        163: new_value_c = 	99;
        164: new_value_c = 	198;
        165: new_value_c = 	145;
        166: new_value_c = 	63;
        167: new_value_c = 	126;
        168: new_value_c = 	252;
        169: new_value_c = 	229;
        170: new_value_c = 	215;
        171: new_value_c = 	179;
        172: new_value_c = 	123;
        173: new_value_c = 	246;
        174: new_value_c = 	241;
        175: new_value_c = 	255;
        176: new_value_c = 	227;
        177: new_value_c = 	219;
        178: new_value_c = 	171;
        179: new_value_c = 	75;
        180: new_value_c = 	150;
        181: new_value_c = 	49;
        182: new_value_c = 	98;
        183: new_value_c = 	196;
        184: new_value_c = 	149;
        185: new_value_c = 	55;
        186: new_value_c = 	110;
        187: new_value_c = 	220;
        188: new_value_c = 	165;
        189: new_value_c = 	87;
        190: new_value_c = 	174;
        191: new_value_c = 	65;
        192: new_value_c = 	130;
        193: new_value_c = 	25;
        194: new_value_c = 	50;
        195: new_value_c = 	100;
        196: new_value_c = 	200;
        197: new_value_c = 	141;
        198: new_value_c = 	7;
        199: new_value_c = 	14;
        200: new_value_c = 	28;
        201: new_value_c = 	56;
        202: new_value_c = 	112;
        203: new_value_c = 	224;
        204: new_value_c = 	221;
        205: new_value_c = 	167;
        206: new_value_c = 	83;
        207: new_value_c = 	166;
        208: new_value_c = 	81;
        209: new_value_c = 	162;
        210: new_value_c = 	89;
        211: new_value_c = 	178;
        212: new_value_c = 	121;
        213: new_value_c = 	242;
        214: new_value_c = 	249;
        215: new_value_c = 	239;
        216: new_value_c = 	195;
        217: new_value_c = 	155;
        218: new_value_c = 	43;
        219: new_value_c = 	86;
        220: new_value_c = 	172;
        221: new_value_c = 	69;
        222: new_value_c = 	138;
        223: new_value_c = 	9;
        224: new_value_c = 	18;
        225: new_value_c = 	36;
        226: new_value_c = 	72;
        227: new_value_c = 	144;
        228: new_value_c = 	61;
        229: new_value_c = 	122;
        230: new_value_c = 	244;
        231: new_value_c = 	245;
        232: new_value_c = 	247;
        233: new_value_c = 	243;
        234: new_value_c = 	251;
        235: new_value_c = 	235;
        236: new_value_c = 	203;
        237: new_value_c = 	139;
        238: new_value_c = 	11;
        239: new_value_c = 	22;
        240: new_value_c = 	44;
        241: new_value_c = 	88;
        242: new_value_c = 	176;
        243: new_value_c = 	125;
        244: new_value_c = 	250;
        245: new_value_c = 	233;
        246: new_value_c = 	207;
        247: new_value_c = 	131;
        248: new_value_c = 	27;
        249: new_value_c = 	54;
        250: new_value_c = 	108;
        251: new_value_c = 	216;
        252: new_value_c = 	173;
        253: new_value_c = 	71;
        254: new_value_c = 	142;
        default: new_value_c = 0;
    endcase
end

always @* begin
    case(alpha_d) //synopsys parallel_case
        0: new_value_d =  1;
        1: new_value_d =  2;
        2: new_value_d =  4;
        3: new_value_d =  8;
        4: new_value_d =  16;
        5: new_value_d =  32;
        6: new_value_d =  64;
        7: new_value_d =  128;
        8: new_value_d =  29;
        9: new_value_d =  58;
        10: new_value_d =  116;
        11: new_value_d =  232;
        12: new_value_d =  205;
        13: new_value_d =  135;
        14: new_value_d =  19;
        15: new_value_d =  38;
        16: new_value_d =  76;
        17: new_value_d =  152;
        18: new_value_d =  45;
        19: new_value_d =  90;
        20: new_value_d =  180;
        21: new_value_d =  117;
        22: new_value_d = 	234;
        23: new_value_d = 	201;
        24: new_value_d = 	143;
        25: new_value_d = 	3;
        26: new_value_d = 	6;
        27: new_value_d = 	12;
        28: new_value_d = 	24;
        29: new_value_d = 	48;
        30: new_value_d = 	96;
        31: new_value_d = 	192;
        32: new_value_d = 	157;
        33: new_value_d = 	39;
        34: new_value_d = 	78;
        35: new_value_d = 	156;
        36: new_value_d = 	37;
        37: new_value_d = 	74;
        38: new_value_d = 	148;
        39: new_value_d = 	53;
        40: new_value_d = 	106;
        41: new_value_d = 	212;
        42: new_value_d = 	181;
        43: new_value_d = 	119;
        44: new_value_d = 	238;
        45: new_value_d = 	193;
        46: new_value_d = 	159;
        47: new_value_d = 	35;
        48: new_value_d = 	70;
        49: new_value_d = 	140;
        50: new_value_d = 	5;
        51: new_value_d = 	10;
        52: new_value_d = 	20;
        53: new_value_d = 	40;
        54: new_value_d = 	80;
        55: new_value_d = 	160;
        56: new_value_d = 	93;
        57: new_value_d = 	186;
        58: new_value_d = 	105;
        59: new_value_d = 	210;
        60: new_value_d = 	185;
        61: new_value_d = 	111;
        62: new_value_d = 	222;
        63: new_value_d = 	161;
        64: new_value_d = 	95;
        65: new_value_d = 	190;
        66: new_value_d = 	97;
        67: new_value_d = 	194;
        68: new_value_d = 	153;
        69: new_value_d = 	47;
        70: new_value_d = 	94;
        71: new_value_d = 	188;
        72: new_value_d = 	101;
        73: new_value_d = 	202;
        74: new_value_d = 	137;
        75: new_value_d = 	15;
        76: new_value_d = 	30;
        77: new_value_d = 	60;
        78: new_value_d = 	120;
        79: new_value_d = 	240;
        80: new_value_d = 	253;
        81: new_value_d = 	231;
        82: new_value_d = 	211;
        83: new_value_d = 	187;
        84: new_value_d = 	107;
        85: new_value_d = 	214;
        86: new_value_d = 	177;
        87: new_value_d = 	127;
        88: new_value_d = 	254;
        89: new_value_d = 	225;
        90: new_value_d = 	223;
        91: new_value_d = 	163;
        92: new_value_d = 	91;
        93: new_value_d = 	182;
        94: new_value_d = 	113;
        95: new_value_d = 	226;
        96: new_value_d = 	217;
        97: new_value_d = 	175;
        98: new_value_d = 	67;
        99: new_value_d = 	134;
        100: new_value_d = 	17;
        101: new_value_d = 	34;
        102: new_value_d = 	68;
        103: new_value_d = 	136;
        104: new_value_d = 	13;
        105: new_value_d = 	26;
        106: new_value_d = 	52;
        107: new_value_d = 	104;
        108: new_value_d = 	208;
        109: new_value_d = 	189;
        110: new_value_d = 	103;
        111: new_value_d = 	206;
        112: new_value_d = 	129;
        113: new_value_d = 	31;
        114: new_value_d = 	62;
        115: new_value_d = 	124;
        116: new_value_d = 	248;
        117: new_value_d = 	237;
        118: new_value_d = 	199;
        119: new_value_d = 	147;
        120: new_value_d = 	59;
        121: new_value_d = 	118;
        122: new_value_d = 	236;
        123: new_value_d = 	197;
        124: new_value_d = 	151;
        125: new_value_d = 	51;
        126: new_value_d = 	102;
        127: new_value_d = 	204;
        128: new_value_d = 	133;
        129: new_value_d = 	23;
        130: new_value_d = 	46;
        131: new_value_d = 	92;
        132: new_value_d = 	184;
        133: new_value_d = 	109;
        134: new_value_d = 	218;
        135: new_value_d = 	169;
        136: new_value_d = 	79;
        137: new_value_d = 	158;
        138: new_value_d = 	33;
        139: new_value_d = 	66;
        140: new_value_d = 	132;
        141: new_value_d = 	21;
        142: new_value_d = 	42;
        143: new_value_d = 	84;
        144: new_value_d = 	168;
        145: new_value_d = 	77;
        146: new_value_d = 	154;
        147: new_value_d = 	41;
        148: new_value_d = 	82;
        149: new_value_d = 	164;
        150: new_value_d = 	85;
        151: new_value_d = 	170;
        152: new_value_d = 	73;
        153: new_value_d = 	146;
        154: new_value_d = 	57;
        155: new_value_d = 	114;
        156: new_value_d = 	228;
        157: new_value_d = 	213;
        158: new_value_d = 	183;
        159: new_value_d = 	115;
        160: new_value_d = 	230;
        161: new_value_d = 	209;
        162: new_value_d = 	191;
        163: new_value_d = 	99;
        164: new_value_d = 	198;
        165: new_value_d = 	145;
        166: new_value_d = 	63;
        167: new_value_d = 	126;
        168: new_value_d = 	252;
        169: new_value_d = 	229;
        170: new_value_d = 	215;
        171: new_value_d = 	179;
        172: new_value_d = 	123;
        173: new_value_d = 	246;
        174: new_value_d = 	241;
        175: new_value_d = 	255;
        176: new_value_d = 	227;
        177: new_value_d = 	219;
        178: new_value_d = 	171;
        179: new_value_d = 	75;
        180: new_value_d = 	150;
        181: new_value_d = 	49;
        182: new_value_d = 	98;
        183: new_value_d = 	196;
        184: new_value_d = 	149;
        185: new_value_d = 	55;
        186: new_value_d = 	110;
        187: new_value_d = 	220;
        188: new_value_d = 	165;
        189: new_value_d = 	87;
        190: new_value_d = 	174;
        191: new_value_d = 	65;
        192: new_value_d = 	130;
        193: new_value_d = 	25;
        194: new_value_d = 	50;
        195: new_value_d = 	100;
        196: new_value_d = 	200;
        197: new_value_d = 	141;
        198: new_value_d = 	7;
        199: new_value_d = 	14;
        200: new_value_d = 	28;
        201: new_value_d = 	56;
        202: new_value_d = 	112;
        203: new_value_d = 	224;
        204: new_value_d = 	221;
        205: new_value_d = 	167;
        206: new_value_d = 	83;
        207: new_value_d = 	166;
        208: new_value_d = 	81;
        209: new_value_d = 	162;
        210: new_value_d = 	89;
        211: new_value_d = 	178;
        212: new_value_d = 	121;
        213: new_value_d = 	242;
        214: new_value_d = 	249;
        215: new_value_d = 	239;
        216: new_value_d = 	195;
        217: new_value_d = 	155;
        218: new_value_d = 	43;
        219: new_value_d = 	86;
        220: new_value_d = 	172;
        221: new_value_d = 	69;
        222: new_value_d = 	138;
        223: new_value_d = 	9;
        224: new_value_d = 	18;
        225: new_value_d = 	36;
        226: new_value_d = 	72;
        227: new_value_d = 	144;
        228: new_value_d = 	61;
        229: new_value_d = 	122;
        230: new_value_d = 	244;
        231: new_value_d = 	245;
        232: new_value_d = 	247;
        233: new_value_d = 	243;
        234: new_value_d = 	251;
        235: new_value_d = 	235;
        236: new_value_d = 	203;
        237: new_value_d = 	139;
        238: new_value_d = 	11;
        239: new_value_d = 	22;
        240: new_value_d = 	44;
        241: new_value_d = 	88;
        242: new_value_d = 	176;
        243: new_value_d = 	125;
        244: new_value_d = 	250;
        245: new_value_d = 	233;
        246: new_value_d = 	207;
        247: new_value_d = 	131;
        248: new_value_d = 	27;
        249: new_value_d = 	54;
        250: new_value_d = 	108;
        251: new_value_d = 	216;
        252: new_value_d = 	173;
        253: new_value_d = 	71;
        254: new_value_d = 	142;
        default: new_value_d = 0;
    endcase
end

always @* begin
    case(value_e) //synopsys parallel_case
        0: new_alpha_e = 0;
        1: new_alpha_e = 0;
        2: new_alpha_e = 1;
        3: new_alpha_e = 25;
        4: new_alpha_e =	2;
        5: new_alpha_e =	50;
        6: new_alpha_e =	26;
        7: new_alpha_e =	198;
        8: new_alpha_e =	3;
        9: new_alpha_e =	223;
        10: new_alpha_e =	51;
        11: new_alpha_e =	238;
        12: new_alpha_e =	27;
        13: new_alpha_e =	104;
        14: new_alpha_e =	199;
        15: new_alpha_e =	75;
        16: new_alpha_e =	4;
        17: new_alpha_e =	100;
        18: new_alpha_e =	224;
        19: new_alpha_e =	14;
        20: new_alpha_e =	52;
        21: new_alpha_e =	141;
        22: new_alpha_e =	239;
        23: new_alpha_e =	129;
        24: new_alpha_e =	28;
        25: new_alpha_e =	193;
        26: new_alpha_e =	105;
        27: new_alpha_e =	248;
        28: new_alpha_e =	200;
        29: new_alpha_e =	8;
        30: new_alpha_e =	76;
        31: new_alpha_e =	113;
        32: new_alpha_e =	5;
        33: new_alpha_e =	138;
        34: new_alpha_e =	101;
        35: new_alpha_e =	47;
        36: new_alpha_e =	225;
        37: new_alpha_e =	36;
        38: new_alpha_e =	15;
        39: new_alpha_e =	33;
        40: new_alpha_e =	53;
        41: new_alpha_e =	147;
        42: new_alpha_e =	142;
        43: new_alpha_e =	218;
        44: new_alpha_e =	240;
        45: new_alpha_e =	18;
        46: new_alpha_e =	130;
        47: new_alpha_e =	69;
        48: new_alpha_e =	29;
        49: new_alpha_e =	181;
        50: new_alpha_e =	194;
        51: new_alpha_e =	125;
        52: new_alpha_e =	106;
        53: new_alpha_e =	39;
        54: new_alpha_e =	249;
        55: new_alpha_e =	185;
        56: new_alpha_e =	201;
        57: new_alpha_e =	154;
        58: new_alpha_e =	9;
        59: new_alpha_e =	120;
        60: new_alpha_e =	77;
        61: new_alpha_e =	228;
        62: new_alpha_e =	114;
        63: new_alpha_e =	166;
        64: new_alpha_e =	6;
        65: new_alpha_e =	191;
        66: new_alpha_e =	139;
        67: new_alpha_e =	98;
        68: new_alpha_e =	102;
        69: new_alpha_e =	221;
        70: new_alpha_e =	48;
        71: new_alpha_e =	253;
        72: new_alpha_e =	226;
        73: new_alpha_e =	152;
        74: new_alpha_e =	37;
        75: new_alpha_e =	179;
        76: new_alpha_e =	16;
        77: new_alpha_e =	145;
        78: new_alpha_e =	34;
        79: new_alpha_e =	136;
        80: new_alpha_e =	54;
        81: new_alpha_e =	208;
        82: new_alpha_e =	148;
        83: new_alpha_e =	206;
        84: new_alpha_e =	143;
        85: new_alpha_e =	150;
        86: new_alpha_e =	219;
        87: new_alpha_e =	189;
        88: new_alpha_e =	241;
        89: new_alpha_e =	210;
        90: new_alpha_e =	19;
        91: new_alpha_e =	92;
        92: new_alpha_e =	131;
        93: new_alpha_e =	56;
        94: new_alpha_e =	70;
        95: new_alpha_e =	64;
        96: new_alpha_e =	30;
        97: new_alpha_e =	66;
        98: new_alpha_e =	182;
        99: new_alpha_e =	163;
        100: new_alpha_e =	195;
        101: new_alpha_e =	72;
        102: new_alpha_e =	126;
        103: new_alpha_e =	110;
        104: new_alpha_e =	107;
        105: new_alpha_e =	58;
        106: new_alpha_e =	40;
        107: new_alpha_e =	84;
        108: new_alpha_e =	250;
        109: new_alpha_e =	133;
        110: new_alpha_e =	186;
        111: new_alpha_e =	61;
        112: new_alpha_e =	202;
        113: new_alpha_e =	94;
        114: new_alpha_e =	155;
        115: new_alpha_e =	159;
        116: new_alpha_e =	10;
        117: new_alpha_e =	21;
        118: new_alpha_e =	121;
        119: new_alpha_e =	43;
        120: new_alpha_e =	78;
        121: new_alpha_e =	212;
        122: new_alpha_e =	229;
        123: new_alpha_e =	172;
        124: new_alpha_e =	115;
        125: new_alpha_e =	243;
        126: new_alpha_e =	167;
        127: new_alpha_e =	87;
        128: new_alpha_e =	7;
        129: new_alpha_e =	112;
        130: new_alpha_e =	192;
        131: new_alpha_e =	247;
        132: new_alpha_e =	140;
        133: new_alpha_e =	128;
        134: new_alpha_e =	99;
        135: new_alpha_e =	13;
        136: new_alpha_e =	103;
        137: new_alpha_e =	74;
        138: new_alpha_e =	222;
        139: new_alpha_e =	237;
        140: new_alpha_e =	49;
        141: new_alpha_e =	197;
        142: new_alpha_e =	254;
        143: new_alpha_e =	24;
        144: new_alpha_e =	227;
        145: new_alpha_e =	165;
        146: new_alpha_e =	153;
        147: new_alpha_e =	119;
        148: new_alpha_e =	38;
        149: new_alpha_e =	184;
        150: new_alpha_e =	180;
        151: new_alpha_e =	124;
        152: new_alpha_e =	17;
        153: new_alpha_e =	68;
        154: new_alpha_e =	146;
        155: new_alpha_e =	217;
        156: new_alpha_e =	35;
        157: new_alpha_e =	32;
        158: new_alpha_e =	137;
        159: new_alpha_e =	46;
        160: new_alpha_e =	55;
        161: new_alpha_e =	63;
        162: new_alpha_e =	209;
        163: new_alpha_e =	91;
        164: new_alpha_e =	149;
        165: new_alpha_e =	188;
        166: new_alpha_e =	207;
        167: new_alpha_e =	205;
        168: new_alpha_e =	144;
        169: new_alpha_e =	135;
        170: new_alpha_e =	151;
        171: new_alpha_e =	178;
        172: new_alpha_e =	220;
        173: new_alpha_e =	252;
        174: new_alpha_e =	190;
        175: new_alpha_e =	97;
        176: new_alpha_e =	242;
        177: new_alpha_e =	86;
        178: new_alpha_e =	211;
        179: new_alpha_e =	171;
        180: new_alpha_e =	20;
        181: new_alpha_e =	42;
        182: new_alpha_e =	93;
        183: new_alpha_e =	158;
        184: new_alpha_e =	132;
        185: new_alpha_e =	60;
        186: new_alpha_e =	57;
        187: new_alpha_e =	83;
        188: new_alpha_e =	71;
        189: new_alpha_e =	109;
        190: new_alpha_e =	65;
        191: new_alpha_e =	162;
        192: new_alpha_e =	31;
        193: new_alpha_e =	45;
        194: new_alpha_e =	67;
        195: new_alpha_e =	216;
        196: new_alpha_e =	183;
        197: new_alpha_e =	123;
        198: new_alpha_e =	164;
        199: new_alpha_e =	118;
        200: new_alpha_e =	196;
        201: new_alpha_e =	23;
        202: new_alpha_e =	73;
        203: new_alpha_e =	236;
        204: new_alpha_e =	127;
        205: new_alpha_e =	12;
        206: new_alpha_e =	111;
        207: new_alpha_e =	246;
        208: new_alpha_e =	108;
        209: new_alpha_e =	161;
        210: new_alpha_e =	59;
        211: new_alpha_e =	82;
        212: new_alpha_e =	41;
        213: new_alpha_e =	157;
        214: new_alpha_e =	85;
        215: new_alpha_e =	170;
        216: new_alpha_e =	251;
        217: new_alpha_e =	96;
        218: new_alpha_e =	134;
        219: new_alpha_e =	177;
        220: new_alpha_e =	187;
        221: new_alpha_e =	204;
        222: new_alpha_e =	62;
        223: new_alpha_e =	90;
        224: new_alpha_e =	203;
        225: new_alpha_e =	89;
        226: new_alpha_e =	95;
        227: new_alpha_e =	176;
        228: new_alpha_e =	156;
        229: new_alpha_e =	169;
        230: new_alpha_e =	160;
        231: new_alpha_e =	81;
        232: new_alpha_e =	11;
        233: new_alpha_e =	245;
        234: new_alpha_e =	22;
        235: new_alpha_e =	235;
        236: new_alpha_e =	122;
        237: new_alpha_e =	117;
        238: new_alpha_e =	44;
        239: new_alpha_e =	215;
        240: new_alpha_e =	79;
        241: new_alpha_e =	174;
        242: new_alpha_e =	213;
        243: new_alpha_e =	233;
        244: new_alpha_e =	230;
        245: new_alpha_e =	231;
        246: new_alpha_e =	173;
        247: new_alpha_e =	232;
        248: new_alpha_e =	116;
        249: new_alpha_e =	214;
        250: new_alpha_e =	244;
        251: new_alpha_e =	234;
        252: new_alpha_e =	168;
        253: new_alpha_e =	80;
        254: new_alpha_e =	88;
        255: new_alpha_e =	175;
        default: new_alpha_e = 0;
    endcase
end

always @* begin
    case(value_f) //synopsys parallel_case
        0: new_alpha_f = 0;
        1: new_alpha_f = 0;
        2: new_alpha_f = 1;
        3: new_alpha_f = 25;
        4: new_alpha_f =	2;
        5: new_alpha_f =	50;
        6: new_alpha_f =	26;
        7: new_alpha_f =	198;
        8: new_alpha_f =	3;
        9: new_alpha_f =	223;
        10: new_alpha_f =	51;
        11: new_alpha_f =	238;
        12: new_alpha_f =	27;
        13: new_alpha_f =	104;
        14: new_alpha_f =	199;
        15: new_alpha_f =	75;
        16: new_alpha_f =	4;
        17: new_alpha_f =	100;
        18: new_alpha_f =	224;
        19: new_alpha_f =	14;
        20: new_alpha_f =	52;
        21: new_alpha_f =	141;
        22: new_alpha_f =	239;
        23: new_alpha_f =	129;
        24: new_alpha_f =	28;
        25: new_alpha_f =	193;
        26: new_alpha_f =	105;
        27: new_alpha_f =	248;
        28: new_alpha_f =	200;
        29: new_alpha_f =	8;
        30: new_alpha_f =	76;
        31: new_alpha_f =	113;
        32: new_alpha_f =	5;
        33: new_alpha_f =	138;
        34: new_alpha_f =	101;
        35: new_alpha_f =	47;
        36: new_alpha_f =	225;
        37: new_alpha_f =	36;
        38: new_alpha_f =	15;
        39: new_alpha_f =	33;
        40: new_alpha_f =	53;
        41: new_alpha_f =	147;
        42: new_alpha_f =	142;
        43: new_alpha_f =	218;
        44: new_alpha_f =	240;
        45: new_alpha_f =	18;
        46: new_alpha_f =	130;
        47: new_alpha_f =	69;
        48: new_alpha_f =	29;
        49: new_alpha_f =	181;
        50: new_alpha_f =	194;
        51: new_alpha_f =	125;
        52: new_alpha_f =	106;
        53: new_alpha_f =	39;
        54: new_alpha_f =	249;
        55: new_alpha_f =	185;
        56: new_alpha_f =	201;
        57: new_alpha_f =	154;
        58: new_alpha_f =	9;
        59: new_alpha_f =	120;
        60: new_alpha_f =	77;
        61: new_alpha_f =	228;
        62: new_alpha_f =	114;
        63: new_alpha_f =	166;
        64: new_alpha_f =	6;
        65: new_alpha_f =	191;
        66: new_alpha_f =	139;
        67: new_alpha_f =	98;
        68: new_alpha_f =	102;
        69: new_alpha_f =	221;
        70: new_alpha_f =	48;
        71: new_alpha_f =	253;
        72: new_alpha_f =	226;
        73: new_alpha_f =	152;
        74: new_alpha_f =	37;
        75: new_alpha_f =	179;
        76: new_alpha_f =	16;
        77: new_alpha_f =	145;
        78: new_alpha_f =	34;
        79: new_alpha_f =	136;
        80: new_alpha_f =	54;
        81: new_alpha_f =	208;
        82: new_alpha_f =	148;
        83: new_alpha_f =	206;
        84: new_alpha_f =	143;
        85: new_alpha_f =	150;
        86: new_alpha_f =	219;
        87: new_alpha_f =	189;
        88: new_alpha_f =	241;
        89: new_alpha_f =	210;
        90: new_alpha_f =	19;
        91: new_alpha_f =	92;
        92: new_alpha_f =	131;
        93: new_alpha_f =	56;
        94: new_alpha_f =	70;
        95: new_alpha_f =	64;
        96: new_alpha_f =	30;
        97: new_alpha_f =	66;
        98: new_alpha_f =	182;
        99: new_alpha_f =	163;
        100: new_alpha_f =	195;
        101: new_alpha_f =	72;
        102: new_alpha_f =	126;
        103: new_alpha_f =	110;
        104: new_alpha_f =	107;
        105: new_alpha_f =	58;
        106: new_alpha_f =	40;
        107: new_alpha_f =	84;
        108: new_alpha_f =	250;
        109: new_alpha_f =	133;
        110: new_alpha_f =	186;
        111: new_alpha_f =	61;
        112: new_alpha_f =	202;
        113: new_alpha_f =	94;
        114: new_alpha_f =	155;
        115: new_alpha_f =	159;
        116: new_alpha_f =	10;
        117: new_alpha_f =	21;
        118: new_alpha_f =	121;
        119: new_alpha_f =	43;
        120: new_alpha_f =	78;
        121: new_alpha_f =	212;
        122: new_alpha_f =	229;
        123: new_alpha_f =	172;
        124: new_alpha_f =	115;
        125: new_alpha_f =	243;
        126: new_alpha_f =	167;
        127: new_alpha_f =	87;
        128: new_alpha_f =	7;
        129: new_alpha_f =	112;
        130: new_alpha_f =	192;
        131: new_alpha_f =	247;
        132: new_alpha_f =	140;
        133: new_alpha_f =	128;
        134: new_alpha_f =	99;
        135: new_alpha_f =	13;
        136: new_alpha_f =	103;
        137: new_alpha_f =	74;
        138: new_alpha_f =	222;
        139: new_alpha_f =	237;
        140: new_alpha_f =	49;
        141: new_alpha_f =	197;
        142: new_alpha_f =	254;
        143: new_alpha_f =	24;
        144: new_alpha_f =	227;
        145: new_alpha_f =	165;
        146: new_alpha_f =	153;
        147: new_alpha_f =	119;
        148: new_alpha_f =	38;
        149: new_alpha_f =	184;
        150: new_alpha_f =	180;
        151: new_alpha_f =	124;
        152: new_alpha_f =	17;
        153: new_alpha_f =	68;
        154: new_alpha_f =	146;
        155: new_alpha_f =	217;
        156: new_alpha_f =	35;
        157: new_alpha_f =	32;
        158: new_alpha_f =	137;
        159: new_alpha_f =	46;
        160: new_alpha_f =	55;
        161: new_alpha_f =	63;
        162: new_alpha_f =	209;
        163: new_alpha_f =	91;
        164: new_alpha_f =	149;
        165: new_alpha_f =	188;
        166: new_alpha_f =	207;
        167: new_alpha_f =	205;
        168: new_alpha_f =	144;
        169: new_alpha_f =	135;
        170: new_alpha_f =	151;
        171: new_alpha_f =	178;
        172: new_alpha_f =	220;
        173: new_alpha_f =	252;
        174: new_alpha_f =	190;
        175: new_alpha_f =	97;
        176: new_alpha_f =	242;
        177: new_alpha_f =	86;
        178: new_alpha_f =	211;
        179: new_alpha_f =	171;
        180: new_alpha_f =	20;
        181: new_alpha_f =	42;
        182: new_alpha_f =	93;
        183: new_alpha_f =	158;
        184: new_alpha_f =	132;
        185: new_alpha_f =	60;
        186: new_alpha_f =	57;
        187: new_alpha_f =	83;
        188: new_alpha_f =	71;
        189: new_alpha_f =	109;
        190: new_alpha_f =	65;
        191: new_alpha_f =	162;
        192: new_alpha_f =	31;
        193: new_alpha_f =	45;
        194: new_alpha_f =	67;
        195: new_alpha_f =	216;
        196: new_alpha_f =	183;
        197: new_alpha_f =	123;
        198: new_alpha_f =	164;
        199: new_alpha_f =	118;
        200: new_alpha_f =	196;
        201: new_alpha_f =	23;
        202: new_alpha_f =	73;
        203: new_alpha_f =	236;
        204: new_alpha_f =	127;
        205: new_alpha_f =	12;
        206: new_alpha_f =	111;
        207: new_alpha_f =	246;
        208: new_alpha_f =	108;
        209: new_alpha_f =	161;
        210: new_alpha_f =	59;
        211: new_alpha_f =	82;
        212: new_alpha_f =	41;
        213: new_alpha_f =	157;
        214: new_alpha_f =	85;
        215: new_alpha_f =	170;
        216: new_alpha_f =	251;
        217: new_alpha_f =	96;
        218: new_alpha_f =	134;
        219: new_alpha_f =	177;
        220: new_alpha_f =	187;
        221: new_alpha_f =	204;
        222: new_alpha_f =	62;
        223: new_alpha_f =	90;
        224: new_alpha_f =	203;
        225: new_alpha_f =	89;
        226: new_alpha_f =	95;
        227: new_alpha_f =	176;
        228: new_alpha_f =	156;
        229: new_alpha_f =	169;
        230: new_alpha_f =	160;
        231: new_alpha_f =	81;
        232: new_alpha_f =	11;
        233: new_alpha_f =	245;
        234: new_alpha_f =	22;
        235: new_alpha_f =	235;
        236: new_alpha_f =	122;
        237: new_alpha_f =	117;
        238: new_alpha_f =	44;
        239: new_alpha_f =	215;
        240: new_alpha_f =	79;
        241: new_alpha_f =	174;
        242: new_alpha_f =	213;
        243: new_alpha_f =	233;
        244: new_alpha_f =	230;
        245: new_alpha_f =	231;
        246: new_alpha_f =	173;
        247: new_alpha_f =	232;
        248: new_alpha_f =	116;
        249: new_alpha_f =	214;
        250: new_alpha_f =	244;
        251: new_alpha_f =	234;
        252: new_alpha_f =	168;
        253: new_alpha_f =	80;
        254: new_alpha_f =	88;
        255: new_alpha_f =	175;
        default: new_alpha_f = 0;
    endcase
end
                   
always @* begin
    case(value_g) //synopsys parallel_case
        0: new_alpha_g = 0;
        1: new_alpha_g = 0;
        2: new_alpha_g = 1;
        3: new_alpha_g = 25;
        4: new_alpha_g =	2;
        5: new_alpha_g =	50;
        6: new_alpha_g =	26;
        7: new_alpha_g =	198;
        8: new_alpha_g =	3;
        9: new_alpha_g =	223;
        10: new_alpha_g =	51;
        11: new_alpha_g =	238;
        12: new_alpha_g =	27;
        13: new_alpha_g =	104;
        14: new_alpha_g =	199;
        15: new_alpha_g =	75;
        16: new_alpha_g =	4;
        17: new_alpha_g =	100;
        18: new_alpha_g =	224;
        19: new_alpha_g =	14;
        20: new_alpha_g =	52;
        21: new_alpha_g =	141;
        22: new_alpha_g =	239;
        23: new_alpha_g =	129;
        24: new_alpha_g =	28;
        25: new_alpha_g =	193;
        26: new_alpha_g =	105;
        27: new_alpha_g =	248;
        28: new_alpha_g =	200;
        29: new_alpha_g =	8;
        30: new_alpha_g =	76;
        31: new_alpha_g =	113;
        32: new_alpha_g =	5;
        33: new_alpha_g =	138;
        34: new_alpha_g =	101;
        35: new_alpha_g =	47;
        36: new_alpha_g =	225;
        37: new_alpha_g =	36;
        38: new_alpha_g =	15;
        39: new_alpha_g =	33;
        40: new_alpha_g =	53;
        41: new_alpha_g =	147;
        42: new_alpha_g =	142;
        43: new_alpha_g =	218;
        44: new_alpha_g =	240;
        45: new_alpha_g =	18;
        46: new_alpha_g =	130;
        47: new_alpha_g =	69;
        48: new_alpha_g =	29;
        49: new_alpha_g =	181;
        50: new_alpha_g =	194;
        51: new_alpha_g =	125;
        52: new_alpha_g =	106;
        53: new_alpha_g =	39;
        54: new_alpha_g =	249;
        55: new_alpha_g =	185;
        56: new_alpha_g =	201;
        57: new_alpha_g =	154;
        58: new_alpha_g =	9;
        59: new_alpha_g =	120;
        60: new_alpha_g =	77;
        61: new_alpha_g =	228;
        62: new_alpha_g =	114;
        63: new_alpha_g =	166;
        64: new_alpha_g =	6;
        65: new_alpha_g =	191;
        66: new_alpha_g =	139;
        67: new_alpha_g =	98;
        68: new_alpha_g =	102;
        69: new_alpha_g =	221;
        70: new_alpha_g =	48;
        71: new_alpha_g =	253;
        72: new_alpha_g =	226;
        73: new_alpha_g =	152;
        74: new_alpha_g =	37;
        75: new_alpha_g =	179;
        76: new_alpha_g =	16;
        77: new_alpha_g =	145;
        78: new_alpha_g =	34;
        79: new_alpha_g =	136;
        80: new_alpha_g =	54;
        81: new_alpha_g =	208;
        82: new_alpha_g =	148;
        83: new_alpha_g =	206;
        84: new_alpha_g =	143;
        85: new_alpha_g =	150;
        86: new_alpha_g =	219;
        87: new_alpha_g =	189;
        88: new_alpha_g =	241;
        89: new_alpha_g =	210;
        90: new_alpha_g =	19;
        91: new_alpha_g =	92;
        92: new_alpha_g =	131;
        93: new_alpha_g =	56;
        94: new_alpha_g =	70;
        95: new_alpha_g =	64;
        96: new_alpha_g =	30;
        97: new_alpha_g =	66;
        98: new_alpha_g =	182;
        99: new_alpha_g =	163;
        100: new_alpha_g =	195;
        101: new_alpha_g =	72;
        102: new_alpha_g =	126;
        103: new_alpha_g =	110;
        104: new_alpha_g =	107;
        105: new_alpha_g =	58;
        106: new_alpha_g =	40;
        107: new_alpha_g =	84;
        108: new_alpha_g =	250;
        109: new_alpha_g =	133;
        110: new_alpha_g =	186;
        111: new_alpha_g =	61;
        112: new_alpha_g =	202;
        113: new_alpha_g =	94;
        114: new_alpha_g =	155;
        115: new_alpha_g =	159;
        116: new_alpha_g =	10;
        117: new_alpha_g =	21;
        118: new_alpha_g =	121;
        119: new_alpha_g =	43;
        120: new_alpha_g =	78;
        121: new_alpha_g =	212;
        122: new_alpha_g =	229;
        123: new_alpha_g =	172;
        124: new_alpha_g =	115;
        125: new_alpha_g =	243;
        126: new_alpha_g =	167;
        127: new_alpha_g =	87;
        128: new_alpha_g =	7;
        129: new_alpha_g =	112;
        130: new_alpha_g =	192;
        131: new_alpha_g =	247;
        132: new_alpha_g =	140;
        133: new_alpha_g =	128;
        134: new_alpha_g =	99;
        135: new_alpha_g =	13;
        136: new_alpha_g =	103;
        137: new_alpha_g =	74;
        138: new_alpha_g =	222;
        139: new_alpha_g =	237;
        140: new_alpha_g =	49;
        141: new_alpha_g =	197;
        142: new_alpha_g =	254;
        143: new_alpha_g =	24;
        144: new_alpha_g =	227;
        145: new_alpha_g =	165;
        146: new_alpha_g =	153;
        147: new_alpha_g =	119;
        148: new_alpha_g =	38;
        149: new_alpha_g =	184;
        150: new_alpha_g =	180;
        151: new_alpha_g =	124;
        152: new_alpha_g =	17;
        153: new_alpha_g =	68;
        154: new_alpha_g =	146;
        155: new_alpha_g =	217;
        156: new_alpha_g =	35;
        157: new_alpha_g =	32;
        158: new_alpha_g =	137;
        159: new_alpha_g =	46;
        160: new_alpha_g =	55;
        161: new_alpha_g =	63;
        162: new_alpha_g =	209;
        163: new_alpha_g =	91;
        164: new_alpha_g =	149;
        165: new_alpha_g =	188;
        166: new_alpha_g =	207;
        167: new_alpha_g =	205;
        168: new_alpha_g =	144;
        169: new_alpha_g =	135;
        170: new_alpha_g =	151;
        171: new_alpha_g =	178;
        172: new_alpha_g =	220;
        173: new_alpha_g =	252;
        174: new_alpha_g =	190;
        175: new_alpha_g =	97;
        176: new_alpha_g =	242;
        177: new_alpha_g =	86;
        178: new_alpha_g =	211;
        179: new_alpha_g =	171;
        180: new_alpha_g =	20;
        181: new_alpha_g =	42;
        182: new_alpha_g =	93;
        183: new_alpha_g =	158;
        184: new_alpha_g =	132;
        185: new_alpha_g =	60;
        186: new_alpha_g =	57;
        187: new_alpha_g =	83;
        188: new_alpha_g =	71;
        189: new_alpha_g =	109;
        190: new_alpha_g =	65;
        191: new_alpha_g =	162;
        192: new_alpha_g =	31;
        193: new_alpha_g =	45;
        194: new_alpha_g =	67;
        195: new_alpha_g =	216;
        196: new_alpha_g =	183;
        197: new_alpha_g =	123;
        198: new_alpha_g =	164;
        199: new_alpha_g =	118;
        200: new_alpha_g =	196;
        201: new_alpha_g =	23;
        202: new_alpha_g =	73;
        203: new_alpha_g =	236;
        204: new_alpha_g =	127;
        205: new_alpha_g =	12;
        206: new_alpha_g =	111;
        207: new_alpha_g =	246;
        208: new_alpha_g =	108;
        209: new_alpha_g =	161;
        210: new_alpha_g =	59;
        211: new_alpha_g =	82;
        212: new_alpha_g =	41;
        213: new_alpha_g =	157;
        214: new_alpha_g =	85;
        215: new_alpha_g =	170;
        216: new_alpha_g =	251;
        217: new_alpha_g =	96;
        218: new_alpha_g =	134;
        219: new_alpha_g =	177;
        220: new_alpha_g =	187;
        221: new_alpha_g =	204;
        222: new_alpha_g =	62;
        223: new_alpha_g =	90;
        224: new_alpha_g =	203;
        225: new_alpha_g =	89;
        226: new_alpha_g =	95;
        227: new_alpha_g =	176;
        228: new_alpha_g =	156;
        229: new_alpha_g =	169;
        230: new_alpha_g =	160;
        231: new_alpha_g =	81;
        232: new_alpha_g =	11;
        233: new_alpha_g =	245;
        234: new_alpha_g =	22;
        235: new_alpha_g =	235;
        236: new_alpha_g =	122;
        237: new_alpha_g =	117;
        238: new_alpha_g =	44;
        239: new_alpha_g =	215;
        240: new_alpha_g =	79;
        241: new_alpha_g =	174;
        242: new_alpha_g =	213;
        243: new_alpha_g =	233;
        244: new_alpha_g =	230;
        245: new_alpha_g =	231;
        246: new_alpha_g =	173;
        247: new_alpha_g =	232;
        248: new_alpha_g =	116;
        249: new_alpha_g =	214;
        250: new_alpha_g =	244;
        251: new_alpha_g =	234;
        252: new_alpha_g =	168;
        253: new_alpha_g =	80;
        254: new_alpha_g =	88;
        255: new_alpha_g =	175;
        default: new_alpha_g = 0;
    endcase
end
        
always @* begin
    case(value_h) //synopsys parallel_case
        0: new_alpha_h = 0;
        1: new_alpha_h = 0;
        2: new_alpha_h = 1;
        3: new_alpha_h = 25;
        4: new_alpha_h =	2;
        5: new_alpha_h =	50;
        6: new_alpha_h =	26;
        7: new_alpha_h =	198;
        8: new_alpha_h =	3;
        9: new_alpha_h =	223;
        10: new_alpha_h =	51;
        11: new_alpha_h =	238;
        12: new_alpha_h =	27;
        13: new_alpha_h =	104;
        14: new_alpha_h =	199;
        15: new_alpha_h =	75;
        16: new_alpha_h =	4;
        17: new_alpha_h =	100;
        18: new_alpha_h =	224;
        19: new_alpha_h =	14;
        20: new_alpha_h =	52;
        21: new_alpha_h =	141;
        22: new_alpha_h =	239;
        23: new_alpha_h =	129;
        24: new_alpha_h =	28;
        25: new_alpha_h =	193;
        26: new_alpha_h =	105;
        27: new_alpha_h =	248;
        28: new_alpha_h =	200;
        29: new_alpha_h =	8;
        30: new_alpha_h =	76;
        31: new_alpha_h =	113;
        32: new_alpha_h =	5;
        33: new_alpha_h =	138;
        34: new_alpha_h =	101;
        35: new_alpha_h =	47;
        36: new_alpha_h =	225;
        37: new_alpha_h =	36;
        38: new_alpha_h =	15;
        39: new_alpha_h =	33;
        40: new_alpha_h =	53;
        41: new_alpha_h =	147;
        42: new_alpha_h =	142;
        43: new_alpha_h =	218;
        44: new_alpha_h =	240;
        45: new_alpha_h =	18;
        46: new_alpha_h =	130;
        47: new_alpha_h =	69;
        48: new_alpha_h =	29;
        49: new_alpha_h =	181;
        50: new_alpha_h =	194;
        51: new_alpha_h =	125;
        52: new_alpha_h =	106;
        53: new_alpha_h =	39;
        54: new_alpha_h =	249;
        55: new_alpha_h =	185;
        56: new_alpha_h =	201;
        57: new_alpha_h =	154;
        58: new_alpha_h =	9;
        59: new_alpha_h =	120;
        60: new_alpha_h =	77;
        61: new_alpha_h =	228;
        62: new_alpha_h =	114;
        63: new_alpha_h =	166;
        64: new_alpha_h =	6;
        65: new_alpha_h =	191;
        66: new_alpha_h =	139;
        67: new_alpha_h =	98;
        68: new_alpha_h =	102;
        69: new_alpha_h =	221;
        70: new_alpha_h =	48;
        71: new_alpha_h =	253;
        72: new_alpha_h =	226;
        73: new_alpha_h =	152;
        74: new_alpha_h =	37;
        75: new_alpha_h =	179;
        76: new_alpha_h =	16;
        77: new_alpha_h =	145;
        78: new_alpha_h =	34;
        79: new_alpha_h =	136;
        80: new_alpha_h =	54;
        81: new_alpha_h =	208;
        82: new_alpha_h =	148;
        83: new_alpha_h =	206;
        84: new_alpha_h =	143;
        85: new_alpha_h =	150;
        86: new_alpha_h =	219;
        87: new_alpha_h =	189;
        88: new_alpha_h =	241;
        89: new_alpha_h =	210;
        90: new_alpha_h =	19;
        91: new_alpha_h =	92;
        92: new_alpha_h =	131;
        93: new_alpha_h =	56;
        94: new_alpha_h =	70;
        95: new_alpha_h =	64;
        96: new_alpha_h =	30;
        97: new_alpha_h =	66;
        98: new_alpha_h =	182;
        99: new_alpha_h =	163;
        100: new_alpha_h =	195;
        101: new_alpha_h =	72;
        102: new_alpha_h =	126;
        103: new_alpha_h =	110;
        104: new_alpha_h =	107;
        105: new_alpha_h =	58;
        106: new_alpha_h =	40;
        107: new_alpha_h =	84;
        108: new_alpha_h =	250;
        109: new_alpha_h =	133;
        110: new_alpha_h =	186;
        111: new_alpha_h =	61;
        112: new_alpha_h =	202;
        113: new_alpha_h =	94;
        114: new_alpha_h =	155;
        115: new_alpha_h =	159;
        116: new_alpha_h =	10;
        117: new_alpha_h =	21;
        118: new_alpha_h =	121;
        119: new_alpha_h =	43;
        120: new_alpha_h =	78;
        121: new_alpha_h =	212;
        122: new_alpha_h =	229;
        123: new_alpha_h =	172;
        124: new_alpha_h =	115;
        125: new_alpha_h =	243;
        126: new_alpha_h =	167;
        127: new_alpha_h =	87;
        128: new_alpha_h =	7;
        129: new_alpha_h =	112;
        130: new_alpha_h =	192;
        131: new_alpha_h =	247;
        132: new_alpha_h =	140;
        133: new_alpha_h =	128;
        134: new_alpha_h =	99;
        135: new_alpha_h =	13;
        136: new_alpha_h =	103;
        137: new_alpha_h =	74;
        138: new_alpha_h =	222;
        139: new_alpha_h =	237;
        140: new_alpha_h =	49;
        141: new_alpha_h =	197;
        142: new_alpha_h =	254;
        143: new_alpha_h =	24;
        144: new_alpha_h =	227;
        145: new_alpha_h =	165;
        146: new_alpha_h =	153;
        147: new_alpha_h =	119;
        148: new_alpha_h =	38;
        149: new_alpha_h =	184;
        150: new_alpha_h =	180;
        151: new_alpha_h =	124;
        152: new_alpha_h =	17;
        153: new_alpha_h =	68;
        154: new_alpha_h =	146;
        155: new_alpha_h =	217;
        156: new_alpha_h =	35;
        157: new_alpha_h =	32;
        158: new_alpha_h =	137;
        159: new_alpha_h =	46;
        160: new_alpha_h =	55;
        161: new_alpha_h =	63;
        162: new_alpha_h =	209;
        163: new_alpha_h =	91;
        164: new_alpha_h =	149;
        165: new_alpha_h =	188;
        166: new_alpha_h =	207;
        167: new_alpha_h =	205;
        168: new_alpha_h =	144;
        169: new_alpha_h =	135;
        170: new_alpha_h =	151;
        171: new_alpha_h =	178;
        172: new_alpha_h =	220;
        173: new_alpha_h =	252;
        174: new_alpha_h =	190;
        175: new_alpha_h =	97;
        176: new_alpha_h =	242;
        177: new_alpha_h =	86;
        178: new_alpha_h =	211;
        179: new_alpha_h =	171;
        180: new_alpha_h =	20;
        181: new_alpha_h =	42;
        182: new_alpha_h =	93;
        183: new_alpha_h =	158;
        184: new_alpha_h =	132;
        185: new_alpha_h =	60;
        186: new_alpha_h =	57;
        187: new_alpha_h =	83;
        188: new_alpha_h =	71;
        189: new_alpha_h =	109;
        190: new_alpha_h =	65;
        191: new_alpha_h =	162;
        192: new_alpha_h =	31;
        193: new_alpha_h =	45;
        194: new_alpha_h =	67;
        195: new_alpha_h =	216;
        196: new_alpha_h =	183;
        197: new_alpha_h =	123;
        198: new_alpha_h =	164;
        199: new_alpha_h =	118;
        200: new_alpha_h =	196;
        201: new_alpha_h =	23;
        202: new_alpha_h =	73;
        203: new_alpha_h =	236;
        204: new_alpha_h =	127;
        205: new_alpha_h =	12;
        206: new_alpha_h =	111;
        207: new_alpha_h =	246;
        208: new_alpha_h =	108;
        209: new_alpha_h =	161;
        210: new_alpha_h =	59;
        211: new_alpha_h =	82;
        212: new_alpha_h =	41;
        213: new_alpha_h =	157;
        214: new_alpha_h =	85;
        215: new_alpha_h =	170;
        216: new_alpha_h =	251;
        217: new_alpha_h =	96;
        218: new_alpha_h =	134;
        219: new_alpha_h =	177;
        220: new_alpha_h =	187;
        221: new_alpha_h =	204;
        222: new_alpha_h =	62;
        223: new_alpha_h =	90;
        224: new_alpha_h =	203;
        225: new_alpha_h =	89;
        226: new_alpha_h =	95;
        227: new_alpha_h =	176;
        228: new_alpha_h =	156;
        229: new_alpha_h =	169;
        230: new_alpha_h =	160;
        231: new_alpha_h =	81;
        232: new_alpha_h =	11;
        233: new_alpha_h =	245;
        234: new_alpha_h =	22;
        235: new_alpha_h =	235;
        236: new_alpha_h =	122;
        237: new_alpha_h =	117;
        238: new_alpha_h =	44;
        239: new_alpha_h =	215;
        240: new_alpha_h =	79;
        241: new_alpha_h =	174;
        242: new_alpha_h =	213;
        243: new_alpha_h =	233;
        244: new_alpha_h =	230;
        245: new_alpha_h =	231;
        246: new_alpha_h =	173;
        247: new_alpha_h =	232;
        248: new_alpha_h =	116;
        249: new_alpha_h =	214;
        250: new_alpha_h =	244;
        251: new_alpha_h =	234;
        252: new_alpha_h =	168;
        253: new_alpha_h =	80;
        254: new_alpha_h =	88;
        255: new_alpha_h =	175;
        default: new_alpha_h = 0;
    endcase
end
endmodule