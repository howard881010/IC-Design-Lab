module test_rop3;

// 1. variable declaration and clock connection
// -----------------------------

// declare variables and connect clock here

// -----------------------------



// 2. connect RTL module 
// -----------------------------

// add your module here

// -----------------------------



// Don't modify this two blocks
// -----------------------------
// input preparation
initial begin
    input_preparation;
end
// output comparision
initial begin
    output_comparison;
end
// -----------------------------


// 3. implement the above two functions in the task file
`include "./rop3.task"


endmodule